`define CPU_CYCLE     1.0 // 100Mhz
`define MAX           800000000 // 3000000
